`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////////////////////////////////////
// Engineer: Abdoula Barry 
// 
// Create Date: 09/27/2024 01:13:00 PM
// Design Name: ArtixNN_digitRecog
// Module Name: digitRecog
// Target Devices: Basys3 Board
// Description: Design of a Digit Finding Neural Network Accelerator using the MNIST Database.
//->Fully parameterized design supporting both ReLU and Sigmoid Activations 
//->Input layer + 4 Layer Design: 784 'input layer' -> 30 layer hidden -> 30 layer hidden -> 10 layer hidden -> 10 layer output
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// AXI4-Lite and AXI Stream Interface
// Using AXI4-Lite and AXI Stream Interface to send unidirectional input data to layer1 of NN
//->More info on AXI found here: https://www.realdigital.org/doc/a9fee931f7a172423e1ba73f66ca4081
/////////////////////////////////////////////////////////////////////////////////////////////////
`include "include.sv"

module digitRecog #(parameter integer C_S_AXI_DATA_WIDTH = 32,
                    parameter integer C_S_AXI_ADDR_WIDTH = 5)
    (
    //Clock and Reset
    input logic s_axi_aclk,
    input logic s_axi_aresetn,
    //AXI Stream Interface - for data to input layer
    input logic [`dataWidth-1:0]            axis_in_data,
    input logic                             axis_in_data_valid,
    input logic                             axis_in_data_ready,
    //AXI Lite Interface
    //->If weights and biases are not configured, the axi lite interface (code generated by IP generator)
    //->allows Processor to communicate with NN
    input logic [C_S_AXI_ADDR_WIDTH-1:0]    s_axi_awaddr,
    input logic [2:0]                       s_axi_awprot,
    input logic                             s_axi_awvalid,
    output logic                            s_axi_awready,
    input logic [C_S_AXI_DATA_WIDTH-1:0]    s_axi_wdata,
    input logic [(C_S_AXI_DATA_WIDTH/8)-1:0] s_axi_wstrb,
    input logic                             s_axi_wvalid,
    output logic                            s_axi_wready,
    output logic [1:0]                      s_axi_bresp,
    output logic                            s_axi_bvalid,
    input logic                             s_axi_bready,
    input logic [C_S_AXI_ADDR_WIDTH-1:0]    s_axi_araddr,
    input logic [2:0]                       s_axi_arprot,
    input logic                             s_axi_arvalid,
    output logic                            s_axi_arready,
    output logic [C_S_AXI_DATA_WIDTH-1:0]   s_axi_rdata,
    output logic [1:0]                      s_axi_rresp,
    output logic                            s_axi_rvalid,
    input logic                             s_axi_rready,
    //Interrupt Interface
    output logic                            intr
    );

    logic [31:0] config_layer_num, config_neuron_num;
    logic [31:0] weightVal, biasVal;
    logic [31:0] out;
    logic out_valid, weightValid, biasValid;

    logic axi_rd_en;
    logic [31:0] axi_rd_data;
    logic softReset;
    
    //for interrupt support so the processor knows when a final output (max value) is found.
    //-> a classification round is finished
    assign intr = out_valid;
    assign axis_in_data_ready = 1'b1;

    //instantiate the axi_lite_wrapper - a customized IP for configuring weights and biases for neurons/links
    axi_lite_wrapper # ( .C_S_AXI_DATA_WIDTH(C_S_AXI_DATA_WIDTH), .C_S_AXI_ADDR_WIDTH(C_S_AXI_ADDR_WIDTH)) 
                    alw (
                        .S_AXI_ACLK(s_axi_aclk), .S_AXI_ARESETN(s_axi_aresetn), .S_AXI_AWADDR(s_axi_awaddr),
                        .S_AXI_AWPROT(s_axi_awprot), .S_AXI_AWVALID(s_axi_awvalid), .S_AXI_AWREADY(s_axi_awready),
                        .S_AXI_WDATA(s_axi_wdata), .S_AXI_WSTRB(s_axi_wstrb), .S_AXI_WVALID(s_axi_wvalid),
                        .S_AXI_WREADY(s_axi_wready), .S_AXI_BRESP(s_axi_bresp), .S_AXI_BVALID(s_axi_bvalid),
                        .S_AXI_BREADY(s_axi_bready), .S_AXI_ARADDR(s_axi_araddr), .S_AXI_ARPROT(s_axi_arprot),
                        .S_AXI_ARVALID(s_axi_arvalid), .S_AXI_ARREADY(s_axi_arready), .S_AXI_RDATA(s_axi_rdata),
                        .S_AXI_RRESP(s_axi_rresp), .S_AXI_RVALID(s_axi_rvalid), .S_AXI_RREADY(s_axi_rready),
                        .layerNumber(config_layer_num), .neuronNumber(config_neuron_num), .weightVal(weightVal),
                        .weightValid(weightValid), .biasValid(biasValid), .biasVal(biasVal),
                        .nnOut_valid(out_valid), .nnOut(out), .axi_rd_en(axi_rd_en),
                        .axi_rd_data(axi_rd_data), .softReset(softReset)
                    );

    logic reset;

    assign reset = ~s_axi_aresetn|softReset;
    // LAYER 1
    //valid signal output from layer1 for each neuron. Technically since all of the neurons will output valid 
    //-> at the same time(due to homogeneous pipelining), only one neurons output can be considered and behavior 
    //-> will remain the same.
    //-> high when neurons have completed activation function execution
    logic [`numNeuronLayer1-1:0] L1_OutValid;
    //L1_TotalOut and L1_HeldDAta represents all the data 'flattened' across every neuron in layer1 for a given activation cycle execution
    logic [`numNeuronLayer1*`dataWidth-1:0] L1_TotalOut, L1_HeldData; 
    logic [`dataWidth-1:0] L1_Out_Data;
    
    layer1 #(.NN(`numNeuronLayer1), .numWeight(`numWeightLayer1), .dataWidth(`dataWidth), .layerNum(1), .sigmoidSize(`sigmoidSize),
             .weightIntWidth(`weightIntWidth), .actType(`Layer1ActType)) 
            L1(
                .clk(s_axi_aclk), .rst(reset), .weightValid(weightValid), .biasValid(biasValid), .weightVal(weightVal),
                .biasVal(biasVal), .config_layer_num(config_layer_num), .config_neuron_num(config_neuron_num), .x_valid(axis_in_data_valid),
                .x_in(axis_in_data), .o_valid(L1_OutValid), .x_out(L1_TotalOut)
            );
    
    //Data from the previous layer is sent serially to all neurons in the next layer by latching the
    //-> full output data to a 'HeldData' register when the layer recieves a valid input signal
    //-> This transfer is implemented using separate FSMs inbetween each layer
    //-> You can imagine a very large shift register inbetween each layer for a hardware representation of the neuron links
    typedef enum {IDLE, SEND} fsm_state;
    fsm_state state_L1SR;
    integer count_1; //counter to represent each neuron; for layer1: counter up to 30 neurons
    logic L1_OutdataValid; //from FSM: send to next layer signaling proper data transfer

    always_ff @(posedge s_axi_aclk) begin
        if(reset) begin
            state_L1SR <= IDLE;
            count_1 <= 0;
            L1_OutdataValid = 1'b0;
        end
        else begin
            case(state_L1SR)
                IDLE: begin
                    count_1 <= 0;
                    L1_OutdataValid <= 1'b0;
                    if(L1_OutValid[0] == 1'b1) begin //neurons have completed execution given an input
                        L1_HeldData <= L1_TotalOut; //Latch the full output data to our held data register
                        state_L1SR <= SEND; //now send the current data
                    end
                end
                SEND: begin
                        L1_Out_Data <= L1_HeldData[`dataWidth-1:0]; //set output data to next layer
                        L1_HeldData <= L1_HeldData >> `dataWidth; //right shift held data to the next data output by our dataWidth
                        count_1 <= count_1+1;//increment count
                        L1_OutdataValid <= 1'b1; //valid data signal to next layer
                        if(count_1 == `numNeuronLayer1) begin //gone through every neuron
                            state_L1SR <= IDLE;
                            L1_OutdataValid <= 1'b0;
                        end
                end
            endcase
        end
    end

    //follow the same convention above for every layer <-to-> layer connection

    // LAYER 2
    logic [`numNeuronLayer2-1:0] L2_OutValid;
    logic [`numNeuronLayer2*`dataWidth-1:0] L2_TotalOut, L2_HeldData; 
    logic [`dataWidth-1:0] L2_Out_Data;
    
    layer2 #(.NN(`numNeuronLayer2), .numWeight(`numWeightLayer2), .dataWidth(`dataWidth), .layerNum(2), .sigmoidSize(`sigmoidSize),
             .weightIntWidth(`weightIntWidth), .actType(`Layer2ActType)) 
            L2(
                .clk(s_axi_aclk), .rst(reset), .weightValid(weightValid), .biasValid(biasValid), .weightVal(weightVal),
                .biasVal(biasVal), .config_layer_num(config_layer_num), .config_neuron_num(config_neuron_num), .x_valid(L1_OutdataValid),
                .x_in(L1_Out_Data), .o_valid(L2_OutValid), .x_out(L2_TotalOut)
            );

    fsm_state state_L2SR;
    integer count_2;
    logic L2_OutdataValid;
    always_ff @(posedge s_axi_aclk) begin
        if(reset) begin
            state_L2SR <= IDLE;
            count_2 <= 0;
            L2_OutdataValid <= 0;
        end
        else begin
            case(state_L2SR)
                    IDLE: begin
                        count_2 <= 0;
                        L2_OutdataValid <= 1'b0;
                        if(L2_OutValid[0] == 1'b1) begin //neurons have completed execution given an input
                            L2_HeldData <= L2_TotalOut; //Latch the full output data to our held data register
                            state_L2SR <= SEND; //now send the current data
                        end
                    end
                    SEND: begin
                            L2_Out_Data <= L2_HeldData[`dataWidth-1:0]; //set output data to next layer
                            L2_HeldData <= L2_HeldData >> `dataWidth; //right shift held data to the next data output by our dataWidth
                            count_2 <= count_2+1;//increment count
                            L2_OutdataValid <= 1'b1; //valid data signal to next layer
                            if(count_2 == `numNeuronLayer2) begin //gone through every neuron
                                state_L2SR <= IDLE;
                                L2_OutdataValid <= 1'b0;
                            end
                    end
            endcase
        end
    end
    
    // LAYER 3
    logic [`numNeuronLayer3-1:0] L3_OutValid;
    logic [`numNeuronLayer3*`dataWidth-1:0] L3_TotalOut, L3_HeldData; 
    logic [`dataWidth-1:0] L3_Out_Data;
    
    layer3 #(.NN(`numNeuronLayer3), .numWeight(`numWeightLayer3), .dataWidth(`dataWidth), .layerNum(3), .sigmoidSize(`sigmoidSize),
             .weightIntWidth(`weightIntWidth), .actType(`Layer3ActType)) 
            L3(
                .clk(s_axi_aclk), .rst(reset), .weightValid(weightValid), .biasValid(biasValid), .weightVal(weightVal),
                .biasVal(biasVal), .config_layer_num(config_layer_num), .config_neuron_num(config_neuron_num), .x_valid(L2_OutdataValid),
                .x_in(L2_Out_Data), .o_valid(L3_OutValid), .x_out(L3_TotalOut)
            );


    //3 LAYER ARCHITECTURE MAXFIND
    logic [`numNeuronLayer3 *`dataWidth-1:0] FinalOutputHeldData;
    assign axi_rd_data = FinalOutputHeldData[`dataWidth-1:0];

    always_ff @(posedge s_axi_aclk) begin
        if(L3_OutValid[0] == 1'b1)  FinalOutputHeldData <= L3_TotalOut;
        else if(axi_rd_en)  FinalOutputHeldData <= FinalOutputHeldData >> `dataWidth;
    end

    //instantiate module to find max output value
    maxFind #(.numInput(`numNeuronLayer3), .inputWidth(`dataWidth))
            MFind(
                .clk(s_axi_aclk), .inData(L3_TotalOut),
                .inValid(L3_OutValid[0]), .outData(out),
                .outValid(out_valid)
            );
endmodule
